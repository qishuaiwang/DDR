
`define DWC_DDRPHY_DFI0_CTRLUPD_ACK_WIDTH 1
`define DWC_DDRPHY_DFI0_CTRLUPD_REQ_WIDTH 1
`define DWC_DDRPHY_DFI0_PHYUPD_ACK_WIDTH 1
`define DWC_DDRPHY_DFI0_PHYUPD_REQ_WIDTH 1
`define DWC_DDRPHY_DFI0_PHYUPD_TYPE_WIDTH 2
`define DWC_DDRPHY_DFI0_DRAM_CLK_DISABLE_WIDTH 1
`define DWC_DDRPHY_DFI0_FREQ_FSP_WIDTH 2
`define DWC_DDRPHY_DFI0_FREQ_RATIO_WIDTH 2
`define DWC_DDRPHY_DFI0_FREQUENCY_WIDTH 5
`define DWC_DDRPHY_DFI0_INIT_COMPLETE_WIDTH 1
`define DWC_DDRPHY_DFI0_INIT_START_WIDTH 1
`define DWC_DDRPHY_DFI0_PHYMSTR_ACK_WIDTH 1
`define DWC_DDRPHY_DFI0_PHYMSTR_CS_STATE_WIDTH 2
`define DWC_DDRPHY_DFI0_PHYMSTR_REQ_WIDTH 1
`define DWC_DDRPHY_DFI0_PHYMSTR_STATE_SEL_WIDTH 1
`define DWC_DDRPHY_DFI0_PHYMSTR_TYPE_WIDTH 2
`define DWC_DDRPHY_DFI0_ADDRESS_WIDTH 6

`define DWC_DDRPHY_DFI0_LP_CTRL_ACK_WIDTH 1
`define DWC_DDRPHY_DFI0_LP_CTRL_REQ_WIDTH 1
`define DWC_DDRPHY_DFI0_LP_CTRL_WAKEUP_WIDTH 5
`define DWC_DDRPHY_DFI0_LP_DATA_ACK_WIDTH 1
`define DWC_DDRPHY_DFI0_LP_DATA_REQ_WIDTH 1
`define DWC_DDRPHY_DFI0_LP_DATA_WAKEUP_WIDTH 5
`define DWC_DDRPHY_DFI0_CTRLMSG_WIDTH 8
`define DWC_DDRPHY_DFI0_CTRLMSG_ACK_WIDTH 1
`define DWC_DDRPHY_DFI0_CTRLMSG_DATA_WIDTH 16
`define DWC_DDRPHY_DFI0_CTRLMSG_REQ_WIDTH 1
`define DWC_DDRPHY_DFI0_ERROR_WIDTH 1
`define DWC_DDRPHY_DFI0_ERROR_INFO_WIDTH 4

`define DWC_DDRPHY_DFI1_CTRLUPD_ACK_WIDTH 1
`define DWC_DDRPHY_DFI1_CTRLUPD_REQ_WIDTH 1
`define DWC_DDRPHY_DFI1_PHYUPD_ACK_WIDTH 1
`define DWC_DDRPHY_DFI1_PHYUPD_REQ_WIDTH 1
`define DWC_DDRPHY_DFI1_PHYUPD_TYPE_WIDTH 2
`define DWC_DDRPHY_DFI1_DRAM_CLK_DISABLE_WIDTH 1
`define DWC_DDRPHY_DFI1_FREQ_FSP_WIDTH 2
`define DWC_DDRPHY_DFI1_FREQ_RATIO_WIDTH 2
`define DWC_DDRPHY_DFI1_FREQUENCY_WIDTH 5
`define DWC_DDRPHY_DFI1_INIT_COMPLETE_WIDTH 1
`define DWC_DDRPHY_DFI1_INIT_START_WIDTH 1
`define DWC_DDRPHY_DFI1_PHYMSTR_ACK_WIDTH 1
`define DWC_DDRPHY_DFI1_PHYMSTR_CS_STATE_WIDTH 2
`define DWC_DDRPHY_DFI1_PHYMSTR_REQ_WIDTH 1
`define DWC_DDRPHY_DFI1_PHYMSTR_STATE_SEL_WIDTH 1
`define DWC_DDRPHY_DFI1_PHYMSTR_TYPE_WIDTH 2
`define DWC_DDRPHY_DFI1_ADDRESS_WIDTH 6

`define DWC_DDRPHY_DFI1_LP_CTRL_ACK_WIDTH 1
`define DWC_DDRPHY_DFI1_LP_CTRL_REQ_WIDTH 1
`define DWC_DDRPHY_DFI1_LP_CTRL_WAKEUP_WIDTH 5
`define DWC_DDRPHY_DFI1_LP_DATA_ACK_WIDTH 1
`define DWC_DDRPHY_DFI1_LP_DATA_REQ_WIDTH 1
`define DWC_DDRPHY_DFI1_LP_DATA_WAKEUP_WIDTH 5
`define DWC_DDRPHY_DFI1_CTRLMSG_WIDTH 8
`define DWC_DDRPHY_DFI1_CTRLMSG_ACK_WIDTH 1
`define DWC_DDRPHY_DFI1_CTRLMSG_DATA_WIDTH 16
`define DWC_DDRPHY_DFI1_CTRLMSG_REQ_WIDTH 1
`define DWC_DDRPHY_DFI1_ERROR_WIDTH 1
`define DWC_DDRPHY_DFI1_ERROR_INFO_WIDTH 4

`include "dfi_prefix_define.sv"

//Customize
`define SVT_DFI_MAX_RANK_WIDTH      `DWC_DDRPHY_DFI0_CS_WIDTH
`define SVT_DFI_MAX_DATA_WIDTH      `DWC_DDRPHY_DFI0_WRDATA_WIDTH
