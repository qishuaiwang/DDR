////////////////////////////////////////
// LPDDR VIP

`timescale 1ps/1fs

`define SVT_LPDDR_MAX_DQ_WIDTH 32

`include "svt_lpddr_full.uvm.pkg"

