`timescale 1ns/1fs
//This module is dummy, used for timescale setting for SDF
`celldefine
module dummy();
endmodule
`endcelldefine
